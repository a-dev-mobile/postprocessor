#######  USER DEFINED EVENTS  #########
##
##     UDE for QTN 200 II MSY and Part Series Technology
##     Andrey V Danilov. St-Petersburg. 24 Apr 2017
##
################################

MACHINE FANUC

#-----------------------------------------------------------------

EVENT qtn_param_take_part
{
   UI_LABEL "MAZAK QTN 200 MSY : Parameters. ������������� : ������ ������."
   CATEGORY MILL DRILL LATHE
   PARAM init_bmp1
   {
      TYPE l
      DEFVAL "${UGII_CAM_USER_DEF_EVENT_DIR}qtn/series_take_part.bmp"
   }

   PARAM qtn_takeover_opt
   {
      TYPE o
      DEFVAL "0. ���������� ����� ���������� #521 #504"
      OPTIONS "0. ���������� ����� ���������� #521 #504","1. ��������� #501 �� ������. #504 ����������.","2. ������������ ������� #501."
      UI_LABEL "����� ������� ���"
   }

   PARAM group_start_1
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "������ ������."
   }
   PARAM qtn_var504
   {
      TYPE s
      DEFVAL "#504"
      TOGGLE Off
      UI_LABEL "����� ������� � ������ ���"
   }
   PARAM qtn_var501
   {
     TYPE d
     DEFVAL "0.0"
     TOGGLE Off
     UI_LABEL "#501 : ���������� ��������� Z2. ����� �� ������"
   }
   PARAM group_end_1
   {
      TYPE g
      DEFVAL "end"
   }

   PARAM group_start_2
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "����. �����. ����."
   }
   PARAM qtn_c2_pos
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "���� ��������� ���"
   }
   PARAM qtn_clrs
   {
      TYPE d
      DEFVAL "1,0"
      TOGGLE Off
      UI_LABEL "���������� �����"
   }
   PARAM qtn_press
   {
      TYPE d
      DEFVAL "0.02"
      TOGGLE Off
      UI_LABEL "������ (�����)"
   }
   PARAM group_end_2
   {
      TYPE g
      DEFVAL "end"
   }

   PARAM group_start_3
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "����������� ����� �������."
   }
   PARAM qtn_var505
   {
      TYPE s
      DEFVAL "#505"
      TOGGLE Off
      UI_LABEL "�������� / ��������� �� / �  ���"
   }
   PARAM qtn_var506
   {
      TYPE s
      DEFVAL "#506"
      TOGGLE Off
      UI_LABEL "����������� �������� ���"
   }
   PARAM group_end_3
   {
      TYPE g
      DEFVAL "end"
   }
}

#-----------------------------------------------------------------

EVENT qtn_param_subspindle_move
{
   UI_LABEL "MAZAK QTN 200 MSY : Parameters. ������������� : �����������"
   CATEGORY MILL DRILL LATHE
   PARAM pull_free_1_expr
   {
      TYPE s
      DEFVAL "#531"
      TOGGLE Off
      UI_LABEL "�������� ��� ������."
   }
   PARAM pull_detal_1_expr
   {
      TYPE s
      DEFVAL "#532"
      TOGGLE Off
      UI_LABEL " �������� � �������."
   }
   PARAM pull_free_2_expr
   {
      TYPE s
      DEFVAL "#533"
      TOGGLE Off
      UI_LABEL "�������� ��� ������."
   }
   PARAM pull_detal_2_expr
   {
      TYPE s
      DEFVAL "#534"
      TOGGLE Off
      UI_LABEL "�������� � �������."
   }
}

#-----------------------------------------------------------------

EVENT qtn_param_subspindle_gohome
{
   UI_LABEL "MAZAK QTN 200 MSY  : Parameters. ����� �������� #2 "
   CATEGORY MILL DRILL LATHE
   PARAM qtn_subspin_gohome_opt
   {
      TYPE o
      DEFVAL "0. ������� ������"
      OPTIONS "0. ������� ������","1. ������� ������","2. �������� � ������� ����������� ������"
      UI_LABEL "����� ������"
   }
   PARAM qtn_var505
   {
      TYPE s
      DEFVAL "#505"
      TOGGLE Off
      UI_LABEL "+ ��������  / - ��������� ���������."
   }
}

#-----------------------------------------------------------------
