#######  USER DEFINED EVENTS  #########
##
##     UDE for QTN 200 II MSY Subspindle
##     Andrey V Danilov. St-Petersburg. 26 apr 2017
##
################################

MACHINE FANUC

#-----------------------------------------------------------------

EVENT qtn_setup
{
   UI_LABEL "MAZAK QTN 200 MSY : ��������� ������"
   CATEGORY MILL DRILL LATHE
   PARAM init_bmp1
   {
      TYPE l
      DEFVAL "${UGII_CAM_USER_DEF_EVENT_DIR}qtn/series_setup.bmp"
   }

   PARAM group_start_1
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "������ ������� ���"
   }
   PARAM qtn_setup_v521
   {
      TYPE d
      DEFVAL "139.0"
      TOGGLE On
      UI_LABEL "#521 : ����� ������� � �������� ���"
   }
   PARAM group_end_1
   {
      TYPE g
      DEFVAL "end"
   }

   PARAM group_start_3
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "������ ������"
   }
   PARAM qtn_setup_var502
   {
     TYPE d
     DEFVAL "50.0"
     TOGGLE Off
     UI_LABEL "#502 : ����� ������� ������"
   }
   PARAM group_end_3
   {
      TYPE g
      DEFVAL "end"
   }
}

#-----------------------------------------------------------------

EVENT barfeeder_list
{
   UI_LABEL "MAZAK QTN 200 MSY : ������ ��� ���������"
   PARAM barfeeder_list
   {
       TYPE   s
       DEFVAL "BARFEEDER_on"
       TOGGLE Off
       UI_LABEL "������ ���������"
   }
}

#-----------------------------------------------------------------

EVENT qtn_subspindle_approach_part
{
   UI_LABEL "MAZAK QTN 200 MSY : ��� : ������ ������."
   CATEGORY MILL DRILL LATHE

   PARAM init_bmp1
   {
      TYPE l
      DEFVAL "${UGII_CAM_USER_DEF_EVENT_DIR}qtn/series_take_part.bmp"
   }

   PARAM group_start_1
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "������ ������"
   }
   PARAM qtn_subspin_takeover_opt
   {
      TYPE o
      DEFVAL "0. ���������� ����� ���������� #521 #504"
      OPTIONS "0. ���������� ����� ���������� #521 #504","1. ��������� �� ������. #504 ����������.","2. ������������ �������� #501."
      UI_LABEL "����� ������� ���"
   }
   PARAM qtn_subspin_v504
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "#504 : ����� ������� � ������ ���"
   }
   PARAM qtn_subspin_v501
   {
     TYPE d
     DEFVAL "0.0"
     TOGGLE Off
     UI_LABEL "#501 : ���������� ��������� Z2. ����� �� ������"
   }
   PARAM group_end_1
   {
      TYPE g
      DEFVAL "end"
   }

   PARAM group_start_2
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "��������� �������"
   }
   PARAM qtn_subspin_c2_pos
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "���� ��������� ���"
   }
   PARAM qtn_subspin_press
   {
      TYPE d
      DEFVAL "0.02"
      TOGGLE Off
      UI_LABEL "������ (�����)"
   }
   PARAM group_end_2
   {
      TYPE g
      DEFVAL "end"
   }

   PARAM group_start_3
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "�������� ����� �������"
   }
   PARAM qtn_subspin_pull
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "�������� / ��������� ������"
   }
   PARAM qtn_subspin_move
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "����������� �������� ���"
   }
   PARAM group_end_3
   {
      TYPE g
      DEFVAL "end"
   }
}

#-----------------------------------------------------------------

EVENT qtn_subspindle_drive
{
   UI_LABEL "MAZAK QTN 200 MSY : ��� : �����������"
   CATEGORY MILL DRILL LATHE

   PARAM init_bmp1
   {
      TYPE l
      DEFVAL "${UGII_CAM_USER_DEF_EVENT_DIR}qtn/move_sub.bmp"
   }
   PARAM init_bmp2
   {
      TYPE l
      DEFVAL "${UGII_CAM_USER_DEF_EVENT_DIR}qtn/move_part.bmp"
   }

   PARAM qtn_move_subspin_1
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "#512 : ����������� ��� ��� ������. +/-"
   }
   PARAM qtn_move_part_1
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "#513 : ����������� ��� � �������. +/-"
   }
   PARAM qtn_move_subspin_2
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "#514 : ����������� ��� ��� ������. +/-"
   }
   PARAM qtn_move_part_2
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "#515 : ����������� ��� � �������. +/-"
   }
}

#-----------------------------------------------------------------

EVENT qtn_subspindle_take
{
   UI_LABEL "MAZAK QTN 200 MSY : ��� : ������� ������ "
   CATEGORY MILL DRILL LATHE
   PARAM qtn_subspin_gohome_opt
   {
      TYPE o
      DEFVAL "0. ������� ������"
      OPTIONS "0. ������� ������","1. ������� ������","2. �������� � ������� ����������� ������"
      UI_LABEL "����� ������"
   }

   PARAM group_start_1
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "������� ������ ���"
   }
   PARAM init_bmp1
   {
      TYPE l
      DEFVAL "${UGII_CAM_USER_DEF_EVENT_DIR}qtn/subspin_free.bmp"
   }
   PARAM qtn_subspin_pull_free
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "#505 : �������� / ��������� ������ �� ���. +/-"
   }
   PARAM group_end_1
   {
      TYPE g
      DEFVAL "end"
   }

   PARAM group_start_2
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "������� ������"
   }
   PARAM init_bmp2
   {
      TYPE l
      DEFVAL "${UGII_CAM_USER_DEF_EVENT_DIR}qtn/subspin_take.bmp"
   }
   PARAM qtn_subspin_move_take
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "#506 : �������� ������� ������� ���. +/-"
   }
   PARAM group_end_2
   {
      TYPE g
      DEFVAL "end"
   }

   PARAM group_start_3
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "�������� ������"
   }
   PARAM init_bmp3
   {
      TYPE l
      DEFVAL "${UGII_CAM_USER_DEF_EVENT_DIR}qtn/subspin_break_off.bmp"
   }
   PARAM qtn_subspin_pull_break
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "#505 : �������� / ��������� ������ �� ���. +/-"
   }
   PARAM qtn_subspin_move_break
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "#506 : �������� ������� ������� ���. +/-"
   }
   PARAM group_end_3
   {
      TYPE g
      DEFVAL "end"
   }
}

#-----------------------------------------------------------------

EVENT qtn_subspindle_m724
{
   UI_LABEL "MAZAK QTN 200 MSY : ��� : �������� ����� �������"
   CATEGORY MILL DRILL LATHE

   PARAM init_bmp1
   {
      TYPE l
      DEFVAL "${UGII_CAM_USER_DEF_EVENT_DIR}qtn/subspin_m724.bmp"
   }
}

#-----------------------------------------------------------------

EVENT qtn_subspindle_cutoff
{
   UI_LABEL "MAZAK QTN 200 MSY : ��� : ������� ���������� ������"
   CATEGORY MILL DRILL LATHE

   PARAM init_bmp1
   {
      TYPE l
      DEFVAL "${UGII_CAM_USER_DEF_EVENT_DIR}qtn/subspin_cutoff.bmp"
   }
}

#-----------------------------------------------------------------
