#######  USER DEFINED EVENTS  #########
##
##     UDE for QTN 200 II MSY
##     Andrey V Danilov. St-Petersburg. 24 Apr 2017
##
################################

MACHINE FANUC

#-----------------------------------------------------------------

EVENT qtn_setup
{
   UI_LABEL "MAZAK QTN 200 MSY : ��������� ������"
   CATEGORY MILL DRILL LATHE
   PARAM init_bmp1
   {
      TYPE l
      DEFVAL "${UGII_CAM_USER_DEF_EVENT_DIR}qtn/series_setup.bmp"
   }

   PARAM group_start_1
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "������ ������� ���"
   }
   PARAM qtn_setup_v521
   {
      TYPE d
      DEFVAL "139.0"
      TOGGLE On
      UI_LABEL "#521 : ����� ������� � �������� ���"
   }
   PARAM group_end_1
   {
      TYPE g
      DEFVAL "end"
   }

   PARAM group_start_3
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "������ ������"
   }
   PARAM qtn_setup_var502
   {
     TYPE d
     DEFVAL "50.0"
     TOGGLE Off
     UI_LABEL "#502 : ����� ������� ������"
   }
   PARAM group_end_3
   {
      TYPE g
      DEFVAL "end"
   }
}

#-----------------------------------------------------------------

EVENT barfeeder_list
{
   UI_LABEL "������ ��� ���������"
   PARAM barfeeder_list
   {
       TYPE   s
       DEFVAL "BARFEEDER_on"
       TOGGLE Off
       UI_LABEL "������ ���������"
   }
}

#---------------------------------------------------------------------------
